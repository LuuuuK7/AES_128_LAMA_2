--	  ________  ________  ________  ___  __    ________  ________  _______           ________  _______   ________      
--	 |\   __  \|\   __  \|\   ____\|\  \|\  \ |\   __  \|\   ____\|\  ___ \         |\   __  \|\  ___ \ |\   ____\     
--	 \ \  \|\  \ \  \|\  \ \  \___|\ \  \/  /|\ \  \|\  \ \  \___|\ \   __/|        \ \  \|\  \ \   __/|\ \  \___|_    
--	  \ \   ____\ \   __  \ \  \    \ \   ___  \ \   __  \ \  \  __\ \  \_|/__       \ \   __  \ \  \_|/_\ \_____  \   
--	   \ \  \___|\ \  \ \  \ \  \____\ \  \\ \  \ \  \ \  \ \  \|\  \ \  \_|\ \       \ \  \ \  \ \  \_|\ \|____|\  \  
--	    \ \__\    \ \__\ \__\ \_______\ \__\\ \__\ \__\ \__\ \_______\ \_______\       \ \__\ \__\ \_______\____\_\  \ 
--	     \|__|     \|__|\|__|\|_______|\|__| \|__|\|__|\|__|\|_______|\|_______|        \|__|\|__|\|_______|\_________\
--	                                                                                                      \|_________|                                                                                                     \|_________|                             
                                                                                                                                          
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use work.my_package.all;

entity rom_invsbox is 

	port (
	clk : in std_logic;
	addr : in std_logic_vector(7 downto 0);
	en   : in std_logic;
	data_out : out std_logic_vector(7 downto 0)
	);
	
end entity;

architecture arch of rom_invsbox is

subtype byte is std_logic_vector (7 downto 0);
  type memory  is array (255 downto 0) of byte;

constant memory_values: memory := (
	 0 => x"52",   1 => x"09",   2 => x"6A",   3 => x"D5",
	 4 => x"30",   5 => x"36",   6 => x"A5",   7 => x"38",
	 8 => x"BF",   9 => x"40",  10 => x"A3",  11 => x"9E",
	 12 => x"81",  13 => x"F3",  14 => x"D7",  15 => x"FB",
	 16 => x"7C",  17 => x"E3",  18 => x"39",  19 => x"82",
	 20 => x"9B",  21 => x"2F",  22 => x"FF",  23 => x"87",
	 24 => x"34",  25 => x"8E",  26 => x"43",  27 => x"44",
	 28 => x"C4",  29 => x"DE",  30 => x"E9",  31 => x"CB",
	 32 => x"54",  33 => x"7B",  34 => x"94",  35 => x"32",
	 36 => x"A6",  37 => x"C2",  38 => x"23",  39 => x"3D",
	 40 => x"EE",  41 => x"4C",  42 => x"95",  43 => x"0B",
	 44 => x"42",  45 => x"FA",  46 => x"C3",  47 => x"4E",
	 48 => x"08",  49 => x"2E",  50 => x"A1",  51 => x"66",
	 52 => x"28",  53 => x"D9",  54 => x"24",  55 => x"B2",
	 56 => x"76",  57 => x"5B",  58 => x"A2",  59 => x"49",
	 60 => x"6D",  61 => x"8B",  62 => x"D1",  63 => x"25",
	 64 => x"72",  65 => x"F8",  66 => x"F6",  67 => x"64",
	 68 => x"86",  69 => x"68",  70 => x"98",  71 => x"16",
	 72 => x"D4",  73 => x"A4",  74 => x"5C",  75 => x"CC",
	 76 => x"5D",  77 => x"65",  78 => x"B6",  79 => x"92",
	 80 => x"6C",  81 => x"70",  82 => x"48",  83 => x"50",
	 84 => x"FD",  85 => x"ED",  86 => x"B9",  87 => x"DA",
	 88 => x"5E",  89 => x"15",  90 => x"46",  91 => x"57",
	 92 => x"A7",  93 => x"8D",  94 => x"9D",  95 => x"84",
	 96 => x"90",  97 => x"D8",  98 => x"AB",  99 => x"00",
	100 => x"8C", 101 => x"BC", 102 => x"D3", 103 => x"0A",
	104 => x"F7", 105 => x"E4", 106 => x"58", 107 => x"05",
	108 => x"B8", 109 => x"B3", 110 => x"45", 111 => x"06",
	112 => x"D0", 113 => x"2C", 114 => x"1E", 115 => x"8F",
	116 => x"CA", 117 => x"3F", 118 => x"0F", 119 => x"02",
	120 => x"C1", 121 => x"AF", 122 => x"BD", 123 => x"03",
	124 => x"01", 125 => x"13", 126 => x"8A", 127 => x"6B",
	128 => x"3A", 129 => x"91", 130 => x"11", 131 => x"41",
	132 => x"4F", 133 => x"67", 134 => x"DC", 135 => x"EA",
	136 => x"97", 137 => x"F2", 138 => x"CF", 139 => x"CE",
	140 => x"F0", 141 => x"B4", 142 => x"E6", 143 => x"73",
	144 => x"96", 145 => x"AC", 146 => x"74", 147 => x"22",
	148 => x"E7", 149 => x"AD", 150 => x"35", 151 => x"85",
	152 => x"E2", 153 => x"F9", 154 => x"37", 155 => x"E8",
	156 => x"1C", 157 => x"75", 158 => x"DF", 159 => x"6E",
	160 => x"47", 161 => x"F1", 162 => x"1A", 163 => x"71",
	164 => x"1D", 165 => x"29", 166 => x"C5", 167 => x"89",
	168 => x"6F", 169 => x"B7", 170 => x"62", 171 => x"0E",
	172 => x"AA", 173 => x"18", 174 => x"BE", 175 => x"1B",
	176 => x"FC", 177 => x"56", 178 => x"3E", 179 => x"4B",
	180 => x"C6", 181 => x"D2", 182 => x"79", 183 => x"20",
	184 => x"9A", 185 => x"DB", 186 => x"C0", 187 => x"FE",
	188 => x"78", 189 => x"CD", 190 => x"5A", 191 => x"F4",
	192 => x"1F", 193 => x"DD", 194 => x"A8", 195 => x"33",
	196 => x"88", 197 => x"07", 198 => x"C7", 199 => x"31",
	200 => x"B1", 201 => x"12", 202 => x"10", 203 => x"59",
	204 => x"27", 205 => x"80", 206 => x"EC", 207 => x"5F",
	208 => x"60", 209 => x"51", 210 => x"7F", 211 => x"A9",
	212 => x"19", 213 => x"B5", 214 => x"4A", 215 => x"0D",
	216 => x"2D", 217 => x"E5", 218 => x"7A", 219 => x"9F",
	220 => x"93", 221 => x"C9", 222 => x"9C", 223 => x"EF",
	224 => x"A0", 225 => x"E0", 226 => x"3B", 227 => x"4D",
	228 => x"AE", 229 => x"2A", 230 => x"F5", 231 => x"B0",
	232 => x"C8", 233 => x"EB", 234 => x"BB", 235 => x"3C",
	236 => x"83", 237 => x"53", 238 => x"99", 239 => x"61",
	240 => x"17", 241 => x"2B", 242 => x"04", 243 => x"7E",
	244 => x"BA", 245 => x"CC", 246 => x"D1", 247 => x"5E",
	248 => x"57", 249 => x"F2", 250 => x"82", 251 => x"47",
	252 => x"AC", 253 => x"E7", 254 => x"2D", 255 => x"95"
	);

begin 
  
  process(clk) is
  begin 
    if rising_edge(clk) and (en = '1') then 
      data_out<= memory_values(to_integer(unsigned(addr)));           
    end if;
  end process;
  
end architecture;